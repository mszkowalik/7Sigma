**$ENCRYPTED_LIB
**$INTERFACE
*$
* TPS43061
*****************************************************************************
* (C) Copyright 2012 Texas Instruments Incorporated. All rights reserved.
*****************************************************************************
** This model is designed as an aid for customers of Texas Instruments.
** TI and its licensors and suppliers make no warranties, either expressed
** or implied, with respect to this model, including the warranties of
** merchantability or fitness for a particular purpose.  The model is
** provided solely on an "as is" basis.  The entire risk as to its quality
** and performance is with the customer
*****************************************************************************
*
* This model is subject to change without notice. Texas Instruments
* Incorporated is not responsible for updating this model.
*
*****************************************************************************
*
** Released by: WEBENCH Design Center, Texas Instruments Inc.
* Part: TPS43061
* Date: 16NOV2012
* Model Type: TRANSIENT
* Simulator: PSPICE
* Simulator Version: 16.2.0.p001
* EVM Order Number: TPS43061EVM-198
* EVM Users Guide: SLVU799November 2012
* Datasheet:
*
* Model Version: Final 1.00
*
*****************************************************************************
*
* Updates:
*
* Final 1.00
* Release to Web.
*
*****************************************************************************
.SUBCKT TPS43061 AGND BOOT COMP EN FB HDRV ISNSN ISNSP LDRV PGND PGOOD
+  PWPD RT_CLK SS SW VCC VIN
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
d054e2d619e668b0706b807646b8037111a8cc64594721807208a85e1aefd30a28587c3a3bc825ce6c6ea971a8291dc76d35d8485846d699639f94b9d14c856a
8f10d309634521e584ae83d57dff2f3582664b04e041863e87b23b8c84a6a67193f17a07f07e954462d766f77596a54b62d6bdea024861df2dd112e4aa362c02
4c365d6473e6054edffda43ce0898750e6479d7d90cea5baf7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
43ff6483192848a26ed53bec7629a4ee165f03a27a1c01fda861090bf3d2be123981d53a6babaa9d3e1786f82095c8a80d71fdea37a778c936361ab795405919
72667800f813325b8dc6150e9752de3228faf8f7a7d9bcd46199f54aea510d32042f0c0c78bb0deb80fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
f197831ab997cb514597b28a3abd988006c017fb2dfda84036806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
2e781867abaac5ce1b1301b16df2da05faa3bfc3f14b9bf72c6ae38325f3cd1495d7fcca0b5012ccddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
2a0dde369b0e03c99162629e90ad3cc673c476259599c8a2278e9f5a89a1ebd0e6b9af996147aa3a589af0812576e61b8318958aa75d4556dd0a70f33e2447ea
4e2689494256295447158635b18b6659ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f62c8b4f8e886a69cc
4b6085f2012636675a0aa31c52cddba976617f42cd5d956bf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
0abb8c42c110d7c51b1301b16df2da051bd7398fd809e6af7e65a63997096a06b032015482838020ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
b0eb42ca922cce59957673035b26e32b2b09d92971e6b7cb6b574213c15e8d89ac5c5dce90c85ba094d295cf8c59dd93473ed35e3f7ec207484379fba1bca2d2
839f52f447781cab957673035b26e32b47d12a5db9c4d228b4bdd1cfb4233b5d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
1e48f80b52cf52581b335ff666912215bd7da830577a40ef1669cf8f0d8f3aa7a873c24146caa13062d6bdea024861df71a419df3b9cd2e17eb34759a160c424
12501895e3f794d935f1882e72da9beadbee2d5133d50126644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
30676e270d7ba14a706b807646b803713c9e038de2490d8707de7db09dabb15462d766f77596a54b62d6bdea024861df71a419df3b9cd2e17eb34759a160c424
b7590adcd9a719c7706b807646b80371467c0f6bb0e0e7b031979312a705a3fd24fdfd9bb2e10b078b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
05146cce2cf93785706b807646b80371c8a933387fb49850ce5ec34e6f8ad1caa5c7c477755fcc9fc0f76534759190ec62d6bdea024861df2dd112e4aa362c02
d9483d90ab4782c2706b807646b80371db78d293143019c49c01dbfd0824bb5b0f090d5b57717962f04163af94c95a1d0d3a4073c77cf9236dc1cba06b961a0c
058bb1d89a84fbf2599bf13f0371d5b42f6ec944424fd010b383949ebd282b37d867a613a0ac2f2b808060ee1504316b5c225826a7752d39aad05fa23ba8b925
6cb87226f48588e51517416927dee8b5ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
179628ee4ab541e880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe2727128158dfa6f6cc90f11a81e844a0bbad8ee659


321c3c0759fb4eb5d6d834f9dcfeac7f29561195cb9a119e2254ae57d4263ab72b3adeaa6c68cb8f8b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
cf260434b9fe12d7706b807646b80371d77001da2bc4ca368492e52ca9907137f9c6ec67082297a00a8cd5950fa7dc893bd627e23244ba5aedfe5c5e91bb342b
317f1bcb1e5ac86291424fe002279da2e1f81912383a31cbf90f7b4f517a06198b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
3b59b36ad64eb58684ae83d57dff2f35a29a80d0fe06482e40aa9f133ccab2462c9ec703c9415b5823b782b3d6a37df173bf76c56446ed39a9a3702383776c53
4c365d6473e6054edffda43ce089875064a66fc0e9ae2280f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
5654d587323d23334a258ad5c6bf4d8a14adece2b524f14cb045613ae43fceace55f5dd8489964f09144f989a85a7e43e384da5d9142d12f2bb0da26e91d20fe
0382627c5bd012d47c3f8de1aca77c883928c3dca9f1370a8c8f7499dfa8f4666606fc3d054efc30c932ea0c66ec2af3a54f0dc4d276ad71b1d22c0c873c0243
1fe70252511a4ce384ae83d57dff2f35b76bbc730b63b4d5bf2c96cea7de6c282cb64a4969cdda32fb39caa823c4ddd76c5cc2503c779cfc5a97c8100a7f5192
66daf9ac6645d3517674bbc8caf0d23de75f53db00dde808838ebe4bcd51da52b34875ad9cf2b042ff7f31d0b5a472a115cde71e5a76569b7928b765497cc849
fe65365436fca01f3fdbae5376dcab6473bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7


5637fcfd860683a9151d9c1419fbf08c7424dd593a343de298f2a95215ae9929693f1203bcc6f135c1cb60b9845d858e24fdfd9bb2e10b072bb0da26e91d20fe
4c365d6473e6054edffda43ce08987500e80a324ba9c4e96f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
4036fe3bb1fccadc151d9c1419fbf08c231ebdeaf0796e4798f2a95215ae9929e8fa70b596afca3f73d9dc50e4e85c45710f626c2faf14a65a97c8100a7f5192
4c365d6473e6054edffda43ce0898750ca391afb5450e0c0f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
2b715364f7d753008dc6150e9752de32af4d796fcbdaa7cbe8c173397f4e2d2624fdfd9bb2e10b078b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
f204860dd3f51380187ea8b1eb3df8de340227790021ef27cea3eb0a2aa7580b5b11621f146daea49a87dce6f28c1cabf04163af94c95a1d58ccff48e3f0f30e
e83d563d614d5ce9d9423b0c849c4a112c3969495f417169b2b0bff6184c43bb24fdfd9bb2e10b078b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
4c365d6473e6054edffda43ce08987503e89331ace5a355fe2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
dbf12f0360092c452fbfcc2b872ff9469e7bf4b828732421ce5ec34e6f8ad1ca5474438ac943e6131652ae74efd59cd45f95a3a83bea06c17612c3486b09b792
7fed2d0d27283289aa33655883cb978b62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b0fb847a3b385fda4597b28a3abd9880fad9ff17a7e9e9d18d0d7d270fe4b7fb6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
b5b551b85673a6bf1b335ff66691221580386cdd3d923a79e8be9181063e91e8cbdebe7801a4e11c41097083f6b3a20980fa21721bf3358cc4169e4a88b5de56
185f27182c5efd10706b807646b80371e76feeb7af3e1b8881a3e6b939a81c4662d766f77596a54b62d6bdea024861df71a419df3b9cd2e17eb34759a160c424
fb1973f283b31bee1b335ff66691221586bdb72f62ea8253677f096f61182f825b11621f146daea49a87dce6f28c1cabf04163af94c95a1d58ccff48e3f0f30e
b64204e7ebac0712c795ec720c2d595e50ba0ae53836ad4c433f2bd729ed5013fbf2872229531c664e462521a6307870a873c24146caa130d7acbf21c6552dd3
4341f824ecf3e2e7706b807646b803719cc4cbb4e93a31fd15b3801d259abfb262d766f77596a54b62d6bdea024861df71a419df3b9cd2e17eb34759a160c424
3e9e5fdcd7dc3d562fbfcc2b872ff94623b96ab753229baa66eaeb9fc4cc8ae16df18951c6eb0f8c474e02c7e8ca851622c8b4d26042e06fd38aff4e12555a5d
256325030bdc7d1e47b82bca135bf5828492e52ca9907137a01a192330666f11f87842ad7aa86c56873aa2fbfbf2d549cb137d57ebc4d10d363b1c9542a67e4a
f18a314737ce6ce36bc5fd38a12d1542ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748


37043a5e33a732b7706b807646b803712e6cec33642d53d10e092ff8d6ec2acbf618abeb8f40b31e710f626c2faf14a66915eb505e8a3b3cfb12c08ee2c37ec0
81bc0cb7c12452441b335ff66691221579e7cd5b00fd645d80d2503a02fcc0716594e2ecfdcb7f1462d6bdea024861df71a419df3b9cd2e17eb34759a160c424
9c3e801b31a04ffe91b0081b127307748415e6c6ba0b32ea6f7fdeb475b80b83077c6957e7dc3aef81951cd64af196171b1caf45b4582faf835b0555b6560412
c3ec163127075deb8dc6150e9752de32c3d5273f1be78e36efea518d467d4be9d37750f413b01fab710f626c2faf14a66915eb505e8a3b3cfb12c08ee2c37ec0
4c365d6473e6054edffda43ce0898750efe11958caf1ca6f8ae76724e38b444f05d79bc20191df12ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
9445347659ec35d3cb3707fed16c224b5a72c2fc6ce7ca51b9a86814d27e1dbd49a56046135d903ded857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
2a76c18f665e8c27be48ce030deefa11ac39e24e6f374294bc41eaf9972019a5aad0cae5ebf3019af04163af94c95a1d0d3a4073c77cf9236dc1cba06b961a0c
0d6a11857a3f7d01f45310c19b6b8ee57e922aa7cbb4b67df88022cc605675ca16767de4da028f5080fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
591d285dfa78c2c64a258ad5c6bf4d8a14adece2b524f14ccb2c584d03eb1e4ca19621dd4ca4acc3c5b57b2266955e82b1d1ca9e44b405a3d7acbf21c6552dd3
8d21fa536185c85c2fbfcc2b872ff9469852c54dc3526c8466eaeb9fc4cc8ae13965adf9533891ac12e89ae99d7349e6aa33655883cb978bd7acbf21c6552dd3
b052355e65d40bda816eb72006c492316867e3e9855280902734814e87d49d0547d9b1cb5fe5d5620fdae27d0c0a851e62d6bdea024861df2dd112e4aa362c02
574f879f1d53d614574ea86a944eba7598f2a95215ae99292652108375a53184fa460eccc75cda6db91f6756c247f62c8b74cc8cf438b7017b9407c104a3fa6d
e72ff3e7fc7190cd07f36db863dd4f4cb162c8e2b10d8623e10bc52e6319ceb0eb9867248335cf44a89afd90dd683fc580fa21721bf3358cc4169e4a88b5de56
d733558f17ca8d9e495b5eae431ecbdcf1e0227cbf3cb102b2bcd6a8bcf625fb13ac6b6121d845c280fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
29fe754104d04f4b706b807646b80371dffa4dce4124f491ce5ec34e6f8ad1ca58ab0039eaebe0d41719d5fa7a267b01ed857e222a29377b9380942fd2fefa16
1f59022967e7ca7b7d49e5986a6ba981d4e4d21d061c186c386b14e28fdab25e12aa4361a7de9e97ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
f594d35fefcc7e2c957673035b26e32b87fe8fb58ba81becb1ca17ffbc42d04873e5642e593a354624fdfd9bb2e10b078b74cc8cf438b7017b9407c104a3fa6d
4c365d6473e6054edffda43ce0898750e339dfcde8e62f5a8ae76724e38b444f05d79bc20191df12ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
3e91d6456c4b63fe706b807646b8037114514c740318c25d2a0eb162ae8d3b98d3b99b01fef3c644a1637079f3d8c51da6b0ac42922a13358ddef45e1d872303
301e882fc7560399ac73e51ea6171029fda4c219b91f031d9d72f8b6ced4c8ae02ad93d405ca8e11ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
658c017bfd47a4cc4597b28a3abd98801d5b620fae8878202c6ae38325f3cd1495d7fcca0b5012ccddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
0360226f8a32fa74e86edc7bbfeb838577292c5f5dee124a212d80903e2d1eaf983b864fed4441a322cff34100050377644126c9831a96bdcad25bf5db12395b
9282ece07efe1537706b807646b803714a213092fd6dee37d960498bee9a6c6c0f090d5b57717962f04163af94c95a1d0d3a4073c77cf9236dc1cba06b961a0c
0fb8138f881bff56706b807646b803717920b9bf903b1b8f118702c88c12390cf418006d7903bf690fa984f27f78bccf9559e1922263399acede045e7c1e1489
3e10a24a415fea9ce027e85c8d068b7373bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
0b00c72b7c2c95cdbe48ce030deefa1195a4122027aef8775a72c2fc6ce7ca5162d7fc06aea0b62b8b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
40ff64b82c572c491aabf11df8bc7d16a1b1eef61449999d8db3ce69c39e6b3543fe2b9debb21178710f626c2faf14a66915eb505e8a3b3cfb12c08ee2c37ec0
4c365d6473e6054edffda43ce089875051095b885b871a6ef7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
a64864cc6ffd637e706b807646b80371610a12217808127f8492e52ca990713707f6b895777902ae82bbfe204ac7c45ee06588b1bf03b89956e2c719886af7e5
014d26bcd4776fef2576175eff3c1c5aed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
3e2f6d3b6fa1f79eddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f63eae6688a631421ee638e7ebcc38d9c4
98b5f0d56fa74586ff1904a7559527c44088a280f80d76dbe10bc52e6319ceb0eb9867248335cf4403a0a7a9237c721380fa21721bf3358cc4169e4a88b5de56
904e90e8e5b2fbfd6ed53bec7629a4ee9cfc4c56529bed119c07274ec8bcb646bafe5040957ee65200d3e0b087c73744ddf7ad811d6a72c444eb3bb0fc4b8a93
4c365d6473e6054edffda43ce0898750daa3a5fb54d4bd36f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
705d459f50f7a08c74114ea99abc715d27be477dbb8da91ab2b0bff6184c43bb24fdfd9bb2e10b078b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
4c365d6473e6054edffda43ce0898750101374417322435ae2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
f637050c6a74cba91b335ff66691221525c511fa5b7513e4138e8d6c9f2df4fc5b11621f146daea49a87dce6f28c1cabf04163af94c95a1d58ccff48e3f0f30e
d5bfd4b79d522d842264a892bdef1efb5d6b58707f577c2f564e1d545515f2e7e9bb8d0e68f5bd5427d9f7e5287cba2c8b74cc8cf438b7017b9407c104a3fa6d
1bd33e665e4e572c6f52d5ca6e23dacf6817b7f0719023cb236e3e8cea9b212773bf76c56446ed39c27a29c2d535fd4ea444f95e85eea42155a6f3f1d348a0ee
abea470061b4cf46495b5eae431ecbdc58207c66a33837180c7b81617ab1e55c2c0fb8a341161179393137f5084e3fa3de4dcf69224b8239ffa02094b80f6ed9
13ac6b6121d845c280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe2727128158dfa6f6cc90f11a81e844a0bbad8ee659
e5e7bd6b4f7f9068706b807646b8037114adece2b524f14c77292c5f5dee124ac1f125687736342ba1d82ae3fd5f9acd00d3e0b087c73744ee626c3c1261d425
4c365d6473e6054edffda43ce08987502d26e210df7c474720b9dfbe3fbec68f96ca58988d555fde73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
59b6ff1c3134b7b51b335ff66691221599a43b8c436cd60d1669cf8f0d8f3aa7a873c24146caa13062d6bdea024861df71a419df3b9cd2e17eb34759a160c424
a22368c484c0be964dec8ad8abd02e9ac1ba77751c81dde0621a54c5698de6ff6969392d5106f0b6a873c24146caa13062d6bdea024861df2dd112e4aa362c02
8807bf206d8a4bf4989c46c74adb5cad9f1fc78125657435a1a90a46f84c8759d16325780afa1b94561ba1e1ffea0410ddf7ad811d6a72c444eb3bb0fc4b8a93
148352bd2f3f1ce3706b807646b8037182218258cca88ffbe7cd59b7f0cb18ab23b782b3d6a37df173bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
8f03dc1d8e018658706b807646b803713ec4349400ec3ee8bd7aac0ae98026628decd1c0ea343a9d6915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
615a28c46d723740bfa54417c4852a036b2e0f7f05f8b6bd55d11f1f786b4406c1cb60b9845d858e24fdfd9bb2e10b078b74cc8cf438b7017b9407c104a3fa6d
4c365d6473e6054edffda43ce08987502bcf036f59aac0c2e2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
94fab6a88c3a1cac74c94f93c383e2571b04712bd5273d12a6908a9fb62203c1042f0c0c78bb0deb80fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
4c365d6473e6054edffda43ce0898750035b8ba07ab513f4f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
94a8023747cab2d9574ea86a944eba7598f2a95215ae9929957be3e376c070904f83950d47b140429c43c24eda4802f7b91f6756c247f62c2bb0da26e91d20fe
abc05a84349f7fe5ac73e51ea6171029fc7da5e9b05a98dbf92a0d9db0bddf19de30493e580a79e6042f0c0c78bb0deb80fa21721bf3358cc4169e4a88b5de56
4c365d6473e6054edffda43ce0898750f8ef2e5cbb06a051e2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
29db0aba6a9e07889551525a7e855e35fee08ee390897965248b8b2b35a0b6c22b3adeaa6c68cb8f8b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
3a31950943f8893e0d0fb41c7f68fd4a1d58caf5355464b56a39eeb6c8f7f3190c7b81617ab1e55cba83e9c74d3a8b7413ac6b6121d845c297636cf94a1578d2
86ad213343ec82a915f60e4ce62d5ce438149ae71d4327b6125916b3dee8ea6e87938bd13c84f8ef042f0c0c78bb0deb80fa21721bf3358cc4169e4a88b5de56
4c365d6473e6054edffda43ce08987501403a0a2c157bd53e2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
1154b5c62790e4722fbfcc2b872ff946b67288f3b0fc30c466eaeb9fc4cc8ae13965adf9533891ac12e89ae99d7349e6aa33655883cb978bd7acbf21c6552dd3
04307dd33841f8905415a1bc588ae6b0449bd2d385565d7f84323401b0599afcd8177ecddd23913c1a23505f6c9c5f8529468a95d6a40ef0a06930635f20c1c3
6c5cc2503c779cfc6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
93d3808648446fd726c880f485e2ca348603798fec049aa28ca9741507fe2e0c00d3e0b087c73744ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
4c365d6473e6054edffda43ce089875055b3f34c08a3b98ae2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
5009e779fac799694dec8ad8abd02e9a2883a51c3334e3143449b260ad47a4b5b032015482838020ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
7142cd1bceb4dc02706b807646b8037134cc3b52a32a1679b2747e3cd181c77e62d766f77596a54b62d6bdea024861df71a419df3b9cd2e17eb34759a160c424
48b4f3abbdab15bb84ae83d57dff2f3500d1d3ebb9c0326796adf5209886a673cb251a2541e3da4c6bc7119ad5724a2a0adedcb26650be7073a3cf9ee36d6dda
1b1caf45b4582faf1b3bd44627b0d1a7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f62c8b4f8e886a69cc
48a94d11d238250fbf139ef5b2461960804b0d8f1855f950a1a90a46f84c8759d16325780afa1b94b270b53054ba30baddf7ad811d6a72c444eb3bb0fc4b8a93
bcd47878fdf46051706b807646b80371ce6505c9fd0ba9d88492e52ca9907137d359fd83916042cd23a80f402716fc46cfaeea42b5578d2f3b300708695416e3
f90824e8f4a0e838706b807646b80371c9790ca48684d169957910123018a02e23b782b3d6a37df173bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
8bf314ab8c034899089653f7e1eda43bf9ca63bb3c278123e10bc52e6319ceb0eb9867248335cf44f5d7409d10e21b7e80fa21721bf3358cc4169e4a88b5de56
f91e9969b8d0883b706b807646b80371be007a8d2a01b1398492e52ca9907137f9c6ec67082297a00a8cd5950fa7dc893ffc32fb7b3a245c3b300708695416e3
6515a1cdba30a506706b807646b803711a96573e18f7381bce5ec34e6f8ad1ca8b415329d984836da92d840fa8f9cb37ed857e222a29377b9380942fd2fefa16
617df87f684e4830a6aef2f846e94004fab5869b49e3f5e1faca85d0862a74fb7e2359a4a403c099e58fadd48448c8c0b4ced54f6781cbe327ab3855428b727c
6d35d8485846d69973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d5f206f4b260aca3e5d0ad1ca54ca84971
b9ed3e04d2a793291b335ff666912215e8fe994e3abed39b33e40e04a931f05f8f22936c7d3b4ad6d3077954e390f95b00d3e0b087c73744ee626c3c1261d425
4c365d6473e6054edffda43ce08987504f64a249ee64d735f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
240cf6a83072ff1a20dd44f77c99c49687647397121a36fa3edf04c157f5dbc073bf76c56446ed39c27a29c2d535fd4ea444f95e85eea42155a6f3f1d348a0ee
c858d814c56a2bccd617b1ae92083d31c9a6d1d11fa70d2e564e1d545515f2e7e9bb8d0e68f5bd547c6a05e67fd634ee8b74cc8cf438b7017b9407c104a3fa6d
6525da4cfd71409daf1922b60cad7ad5a40b0129de2089fb62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a96f3b666d9ed3040f
81a9746d786d11d6151d9c1419fbf08ca96da287e296fcafd392b39ab991fc45be65b7c13d451c0d12aa4361a7de9e97b03201548283802070870f25f43711dd
c8ec67115e15a9b2ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f63eae6688a631421ee638e7ebcc38d9c4
09f36a1d8b68f4d8151d9c1419fbf08ce6d075e2ee7e9a255a444ae3de1b9453977aa12e8ea1263dbaa78b47fb353ab3f04163af94c95a1d58ccff48e3f0f30e
c0ff0c48b49f7f3384ae83d57dff2f3528465d875bdfcfd798f2a95215ae9929ae81c35cd84c1fbb49bcb2e9b7241eb4644126c9831a96bdcad25bf5db12395b
4c365d6473e6054edffda43ce0898750dcdf8d7f3c517bc8f7869ff373847bc78cb450af0c5bc3638b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
b0686e6017586587706b807646b803714aa29e307ae1bf81ce5ec34e6f8ad1caa5c7c477755fcc9f4d65a3db4bba07aaed857e222a29377b9380942fd2fefa16
5ff44a992c4e2ee34597b28a3abd9880c4e73f9938a3cefc7e65a63997096a06b032015482838020ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
62748d827ca277c7706b807646b80371c83805c2174809e866eaeb9fc4cc8ae10d84fbc6657014080b4a1f9401332bc16d35d8485846d699639f94b9d14c856a
58ab99932615660b1b335ff666912215c05799f034d3e1609bb32ef3089dcfcfdad4b7980b83d60c73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
04f5acd939422ec02dce7963c39dbc2ecdbcb8ac08cc1915faca85d0862a74fbceff41e4364046085e09e353ec4d4fa516e3ac88ef572561e84db9cc2173f1ad
8a974bc2a1288303ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
0805c9bc4a8c6e82b9d15c5be4e02d4923d50fbd82f4809ad8d46728fbe449b87cc7b74c860f658f67138a307a6c221bb91f6756c247f62c2bb0da26e91d20fe
8c74ba1df3e17c1c706b807646b803718d9d46dab323e282a09546df2e73c22f7236390f27aa280755bd0a8bf739c7dece523d51c4bd91cd2bb0da26e91d20fe
d36d26370afc449b1b1301b16df2da0573d332867f5790aced857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
394197bedeb77a71d05ee9f4a2babc05a378d1a54122e7f1bde2f9726e2f693dff3863bf4c9cdd7724fdfd9bb2e10b078b74cc8cf438b7017b9407c104a3fa6d
4c365d6473e6054edffda43ce08987508c655ab34a33bf3fe2ba4357ad2ad1ff421e1c7e544985036915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
0309faec1d3e3fba706b807646b80371da0990a7c75136fd187a22d5c7ce302bfaeaa281e22d723e644126c9831a96bdf04163af94c95a1d58ccff48e3f0f30e
47e2519fa42d321e84ae83d57dff2f3522b88249def5964b96adf5209886a673a027d9bf4111f52d2d3711465512234c9a87dce6f28c1cabcad25bf5db12395b
b9ac294d39eede85187ea8b1eb3df8de4a96d889436bba3ba6db312667ee6b9fa873c24146caa13062d6bdea024861df71a419df3b9cd2e17eb34759a160c424
d8d4f554fe5763de29e825b94f56ec70eaddf1740b36e06fa1b8e96d36cb7a52dad4b7980b83d60c73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
53428b3d5fabd5e9706b807646b80371b2a722aeccdc78b9ef444a8a0e181a19f618abeb8f40b31e710f626c2faf14a66915eb505e8a3b3cfb12c08ee2c37ec0
ab826d58a5e292c658e7dc8c8e0923333fe71322b6154693726d9a7f6b37359c1b3bd44627b0d1a7ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
30121bf0e4b6f88026c880f485e2ca34c7ae5a91fde77d89e5ff990aaf2cc607ed857e222a29377b14aee5f82b16b7673d4db86b42817e2bf411d12d7ec6c2f4
c9df73872fc60450fe4e3ad5ef653a2c64cb1cfefb6e4006017f6156319502eb86dfd129f9d4d35e826d63767c184704644126c9831a96bdcad25bf5db12395b
19783a1fc48c2a0c78ffbc956a033e59506f70b030c78a07019b8717068e3d44e10bc52e6319ceb0eb9867248335cf444b1ed20257b6422a639f94b9d14c856a
f80a395284a571112fbfcc2b872ff94650d47cfb7ccb7fdb66eaeb9fc4cc8ae13965adf9533891ac030135283f2f4fe7b0655b7297d2cc5b1aabfa10941d45cf
f9705fba3e9419e84a749c3c8ff77c97ecd04b518e08577bf6b416f84d54d658844da759261db9866915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
e080b6f7611af9f11b335ff666912215eddb52431de15019a00c9e422d3f61ec8a839d41e6673fceb58626e19d95465c3b2051e815b1bd147a800e49a4c57238
c2c5719688b9adbb62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b581739c5c1ab2d23f214b807900fe3ac5c
099a86bb88e9bfe3495b5eae431ecbdce1e890e7986dcba2d18e72a97ccdabb1fb39caa823c4ddd76c5cc2503c779cfc6915eb505e8a3b3cfb12c08ee2c37ec0
e9dd452c4e6cfebe969deb1afc4fde25764eb50ebf3f76adf79ed346fe02bf5df04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
fe9073afece57ff8706b807646b803718ea1fd7daa70489b8492e52ca9907137f9c6ec67082297a00a8cd5950fa7dc899542b05b8572c0993b300708695416e3
a2bf575280f8d8aaf45310c19b6b8ee5e8be9181063e91e8d565d3fae6b810699c43c24eda4802f7b91f6756c247f62c8b74cc8cf438b7017b9407c104a3fa6d
4559754b57dd997c42267015cdc870b232b6d9b65cadb3c02c6ae38325f3cd1495d7fcca0b5012ccddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
efaf3b99682e31791b335ff666912215fb6f1944dc560567825288324a0dbaed1c64e4fae4013ac4e41f235217d54a8da5dd93e2580e537f639f94b9d14c856a
52ba738fba12eb4af959dbdbcb8ecc1be7c9776c786c195880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
a61e1bc8f3d9b1db26c880f485e2ca34c337c4bc72c91cb47870b400afe279c562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
881857014bf756d4706b807646b8037187e4345caa5828648492e52ca99071370f644d38cd9290e17582c6bfc3c5e874fe5fca639a680f688ddef45e1d872303
e6573f93da02bfe7b66f5818b430d8dcd3f5f1cb4e78ae962c6ae38325f3cd1495d7fcca0b5012ccddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
2215305de2bb21fe151d9c1419fbf08c255a9f07e5655ff27d4e8ec01023cbc998f2a95215ae9929589af0812576e61b1b3bd44627b0d1a7ee626c3c1261d425
846dad09021724e51b335ff666912215af4c491e4418dbeaa0c624c3e799bda573bf76c56446ed39c27a29c2d535fd4ea444f95e85eea42155a6f3f1d348a0ee
a9174ed1bf108f9a4f83950d47b14042446e981d06afb3c5ab9e97ff8c1f9167e55f5dd8489964f09144f989a85a7e43c612182fe29e690d5a97c8100a7f5192
96a13383adcb4a430d0fb41c7f68fd4a82c3f834928beb5e553d7b0be28304d5726d9a7f6b37359c1b3bd44627b0d1a7ddf7ad811d6a72c444eb3bb0fc4b8a93
0e93a9674d9c6bf6706b807646b8037152640ce34dd7f4088492e52ca9907137a01a192330666f11e7349691d690240f72a4cd21040a3877ea3882c684659db1
224fe9df4b4ef4f2b9d15c5be4e02d49b25b708b842430b7726d9a7f6b37359c1b3bd44627b0d1a7ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
1333f3c86417d3f201e07779432d240b7be5161367a34e4c6b574213c15e8d895f22b35d16ee0ba8b3715af44a0e252df44496155f03ed4fd7acbf21c6552dd3
$CDNENCFINISH
.ENDS TPS43061
*$
.subckt TPS43061_TOPLEVEL_S10 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
2c5ce0287ce5ddeb46b92e86e8aaa0ba77968c367c5eb47975ba0c3b03da98f26915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
39deafbe7a97ca4d1852d2bae25628728884162488a3797780fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
1e7e75f62a07f7b1bbcb463bf6330e44495a9bb7954552cde75adc0303e81669422d94caab3a0e7ed9341a119a21aaf1b4a02f072722f4b52cf859073b56ae0f
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S10
*$
.subckt TPS43061_TOPLEVEL_S11 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
e78fee54ef52378d46b92e86e8aaa0ba77968c367c5eb479879f0c9fbb8e40016915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
699fd6531918f3dc1852d2bae25628728884162488a3797780fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
1e7e75f62a07f7b1bbcb463bf6330e44575ba129fd85412be75adc0303e81669beac70612beb6e179ea5842bf7c428edb4a02f072722f4b52cf859073b56ae0f
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S11
*$
.subckt TPS43061_TOPLEVEL_S2 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
c21144fd15b2c61331820e631d1d1d7423f284e2e346bfb8ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
e07b7a6acd4bf43c6f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44eff574bcdcb677aa0ffb76e2ddf4497b2b7447af30eda7a9af673fe4a4241386e23b0d90c7c299fe6e2969c0b1ba3f40
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S2
*$
.subckt TPS43061_TOPLEVEL_S5 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
a41eff5afcadbe0431820e631d1d1d74cce714c3daebb9efed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
0d00147a4ec8159a6f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e444ffca53f33c7306d0ffb76e2ddf4497b2b7447af30eda7a94581845dadf41c9e1af09922ee8b758c1170ec9fe77f9354
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S5
*$
.subckt TPS43061_TOPLEVEL_S12 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
a2bb1bfa319d55b546b92e86e8aaa0ba77968c367c5eb4792f2bd09e50f291d26915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
eef19482dea315b11852d2bae25628728884162488a3797780fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
1e7e75f62a07f7b1bbcb463bf6330e445c12dbc36bfd1b6ae75adc0303e81669beac70612beb6e175fbb6ccbaa4bb091e23b0d90c7c299fe6e2969c0b1ba3f40
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S12
*$
.subckt TPS43061_TOPLEVEL_S3 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
49437a5c2c000e5531820e631d1d1d7451c16968e1146dc5ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
196545b3a77859896f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e449fca2d09a1602b870ffb76e2ddf4497b2b7447af30eda7a9fe99c2387d62d51db4a02f072722f4b52cf859073b56ae0f
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S3
*$
.subckt TPS43061_TOPLEVEL_S6 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
984f32a07473fb7c31820e631d1d1d74ef1e214e65ee9ca6ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
dd1eb1f7fd6960a06f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44dd4a5f3ed5996b330ffb76e2ddf4497be9ba6df74be059f8e421b088f586f07d1af09922ee8b758c1170ec9fe77f9354
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S6
*$
.subckt TPS43061_TOPLEVEL_S7 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
ca116cfd9f503f5a31820e631d1d1d74bc43870b2068c893ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
22fa704315324fee6f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44b8257e7c370c44b80ffb76e2ddf4497b2b7447af30eda7a94581845dadf41c9e1af09922ee8b758c1170ec9fe77f9354
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S7
*$
.subckt TPS43061_TOPLEVEL_S1 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
44f117741689d59131820e631d1d1d749e35700c7913e939ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
3c76beba9b808c126f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e447b3ba2fd65dbf9050ffb76e2ddf4497b2b7447af30eda7a926c4639be54aeef78ed77f303759ed3ce236655da4ddb080
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S1
*$
.subckt TPS43061_TOPLEVEL_S8 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
48cad54cbc66f42d31820e631d1d1d740e2409c315f54deced857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
e65d04c3f5d7c4236f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44a0cccacb04419cb30ffb76e2ddf4497be9ba6df74be059f8e421b088f586f07d1af09922ee8b758c1170ec9fe77f9354
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S8
*$
.subckt TPS43061_TOPLEVEL_S4 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
cca5ca7cd3bb954631820e631d1d1d743397604f987b60beed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
c89815736fd06a736f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44d3c3547c91af769e0ffb76e2ddf4497b2b7447af30eda7a917bce6db3835e7a3e23b0d90c7c299fe6e2969c0b1ba3f40
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S4
*$
.subckt TPS43061_TOPLEVEL_F1 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
ae601cf82fbefc0c31820e631d1d1d74872d6da6e74e75eeed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
969b68e4450fa8bd6f31076d2b37e96b3a7bc5327c69eeafddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_F1
*$
.subckt TPS43061_TOPLEVEL_S13 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
cac64a474f6db0d746b92e86e8aaa0ba77968c367c5eb479ed483728f87a2ff56915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
204d864dd5c51c161852d2bae25628728884162488a3797780fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
1e7e75f62a07f7b1bbcb463bf6330e442a2f0d2b46524d4ce75adc0303e81669cb43e85d9037ba9df9bca68dcba27aa0a199dc71632da75a15fea89cf14f6bad
595b7ea07c82f5178b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S13
*$
.subckt TPS43061_TOPLEVEL_S9 1 2 3 4
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
0d4fba81348870d631820e631d1d1d74525a947d4222b598ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
7e9baaa9719bd1f96f31076d2b37e96baa35006d782c6ce9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1e7e75f62a07f7b1bbcb463bf6330e44ccbbb1088960694e0ffb76e2ddf4497b2b7447af30eda7a926c4639be54aeef7c86660c3d13115677ab4b31efee64103
$CDNENCFINISH
.ends TPS43061_TOPLEVEL_S9
*$


** Wrapper definitions for AA legacy support **


.subckt d_d1 1 2


$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
1580a2664af5c9b71dffb53947c4a0506915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f


0697746efb67a3a341e6e617f9adb744ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f62c8b4f8e886a69cc
f7a854a98d732f8b65b706867a9136e68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
39c84b0c9f72e0078e024cbd033ee0af8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
0660a0f5c4a1d536aad0cae5ebf3019af04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
eff9bf1926aa5ce162d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b581739c5c1ab2d23f214b807900fe3ac5c


$CDNENCFINISH
.ends d_d1


.subckt d_d 1 2


$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
1580a2664af5c9b79ba351c972f8011bf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb


0697746efb67a3a37eef396dcc27bc378b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
f7a854a98d732f8b65b706867a9136e68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
017be23040227359ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
39c84b0c9f72e0078e024cbd033ee0af8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941


$CDNENCFINISH
.ends d_d


*$
.SUBCKT csd86330q3d  1 2 3 4 5 6 7 8 9
*
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
7dc8e005cc47bb4dfd56be15e936ee27236003f871c85c940a746c3bc2d639d88b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
0c4550fdccd06d4af4305df9f983f209f1d13c678e4e9d7b3f1d1223929dfd898b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
2eab0b400fa84ed703aa89060feebfaa55eec14a850e369ebe4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
5505adfa69bc3d25319cc27e7cf4b89a17c31722fb1fdba8be4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
d2d6a088b20ade6d9aac079c398971b9854178155f52c3968cd0517f0151e5d08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
b3f21c82fe924a3e7f28d33e21cfb73a854178155f52c3968cd0517f0151e5d08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
a533432b48c3a0cc87d80f094815c07755eec14a850e369ebe4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
84e3b35d4c9fdb652f1eb6baad5d55e9651630069b2345f46e1558c1d8d21db5ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
9496bdcf840f5f77d58aa4bf425b181d651630069b2345f46e1558c1d8d21db5ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
0d9cc6e38e7abb6311d8cb30cfa55420651630069b2345f46e1558c1d8d21db5ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
544704b4c918a8072db3696be623eff76c11c24ae712f9afc1a23a0a43bd134480fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd5469306ad371de54
91efe665173dc491608158c389b4ff3f0668b7fba1edb69efc38f1d98ada2dc9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
50522329b8a8b20813f02cc56ee30f07651630069b2345f424a28f27ab473008ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
c3abad7d0bf5ffc92c7834446899169b121475774a964e71ddd213233cbbfb79ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
6fe68377a0ae8f902c7834446899169bf02523f77385cf5c73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
ce87a7d05ebe4457fafa402b4ddf25c90668b7fba1edb69efc38f1d98ada2dc9ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
701bb725b19e8ea871375c2e82ac9b18bf6602dce5bbf22dddd213233cbbfb79ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
$CDNENCFINISH
.ENDS csd86330q3d
**********************************************************************
**********************************************************************
*                                                                    *
*   n36306   -  PSpice Model                                         *
*                                                                    *
*   n36306 is the LS silicon die model for use with 86330q3d         *
*                                                                    *
**********************************************************************
**********************************************************************
* SUBCKT Definition:  1=D  2=G  3=S
**********************************************************************
.SUBCKT n36306  1 2 3
* PARAMETER (local) DEFINITIONS SECTION
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
2cfd781695004e385100148e3d6e300dd7ca745dc7133bfb62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a96f3b666d9ed3040f
2cfd781695004e387bc7ce494a63b95cab4f8f49c9687b8980fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
2cfd781695004e38126b113ea1f9ad80423ac9b346247ddb60c5ac4de13f4064ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
2cfd781695004e383edbcd936276c8ebc5329e5ca5bcd06519842dc9a1099cd50399937abc26ad30c3444eda896b7868ed857e222a29377b9380942fd2fefa16
2cfd781695004e38444ffe5a14ddde1869dc209837ee3cb473bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
****** MODEL SUBCIRCUIT BEGINS HERE     ******************************
1387a7647ddaf4b444ba8c84c92e471c90b8469c307059f0743db0b1d721bf3b93e9a193d756852ed0afb64e782c9040d6123d4363d6790fb2a0eb8b33b5b074
bb2d40765b665fa96915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
d3ae90bb1cd66be0e04afeef43cc7d7162d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
cbe37d5098e0c17857e7d96e6be9ec93d76bf3d4fbc8a367ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
6401eb28bd845c08b1fface195ae7535ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
f569dfd879b574769bf727f497549dda39859341766fc92cf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
7a13c2b4abc7a0c32a73071912eabad1ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
1bf2775e5d19f4618255cd4c1295482d39859341766fc92cf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
35a1ca33872f2041c6619b7646f07228049104bb5d4ca56dbe401a404cd83ba166fa3ae85270d163ea2cf4e7d413dba4c2ec0d54e1fbf00c21ee64457ea555af
13daf902c18c20b08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
5547dc123c3fce4b4c6e15a319498476c7541ec212b25801f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
3ebc5ddc64c3d282562cd66acf34399062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b324271c0280911f7df87e9386ba9e8f62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
22118ccc9a4693cb403ec2eb20ef56aced857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
5b8be7694daebfb6b95dbd4ca0a9140c3e97f995c31a36e776617f42cd5d956bf04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
15aa5a803ed33c3095e6484c921cd1d92d973a8ca393d7ffbe4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
5cc23a905735a528a38cbb9f2df12dda063cd1b01c757500be4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
*******************************************************************
1e7e75f62a07f7b186e471729bc5541749b5e96410c30f2547f3e73fa04e71d0c24394b0aefd2664706b807646b80371ba80e3b7e443da4b4f85a241c9207b84
262b99977648e9d16c5e49ef621538cd706b807646b80371d3a99143ac7ecc477696203bced13e84f80c4c8e2b766bd8824901d9f53d509df4c83cab6b9aced6
b27e2e819491226c0e8f570a764b71b1b61718b66f0797759c23c515e4041152361bb2002e6a78c008e79cbf8de54de39a283b42b20f2dfbef2b9269f316b7f3
809d1592585346e42410f9b01f28bfc2706b807646b80371401e692c311d9e41fe670db4bdff8f92706b807646b80371c3be9dd39875721b6b8f064b73f0f573
a284042cd791aa6e878b30bcf251304b706b807646b80371ea35a63cd16a7017fe670db4bdff8f92706b807646b803718c2889ca49ca0fe3d0a7caf6cdbb631c
3b1feb6bf520a7922c91fded96c93703f6a2b547dc976ba0bb29955bae8f226f4005379e431e12f3b585b96681e0ca9bfe3ce9cf33d8558c68957789b47fb3f9
4134e00fa366ca83e238000989aa4a17f6a2b547dc976ba039b302d18fa67a4265e99d0d47459603a84ecbc7159c51adad084f03a18c1696f62496a6a101fce4
9e13f6a7b30c0d5837ae7c67df5f62a1706b807646b8037134c64911cb9a3b9ae3568e8b165a35ba706b807646b8037128b2f6472235ee1ed9cd054cffe4113f
a6b5fbf4542e095a6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
7b0faa21729cd1dcc65fa3fd5d6e3745706b807646b80371e84c4e9059d274e77a74c1a9b086f5a93421bf8d63a79fc975ae2546e9b9532925bae6d262f7a4f8
5f57011c64ecdeb2e30dea4b4d29e81b706b807646b80371d01a699e884848be787f0235f323548f706b807646b80371c5ed5780386810ae655e130736f46d73
41076da6468fadded813ef29de50e822706b807646b80371e80dcfcbc57bfea86f0b6265b9122619706b807646b803718b03d7c2720630032e80e42bd2ee1bc1
03dc106fabbcecab6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
f8877d765eca4de053e46a310f19d695706b807646b803712b20e00307d47b5ecdf9f7c3abc57dae706b807646b80371bb98c84c0bea3b3eb4537737a844a535
1b56e1e057d96a20135c898b90113bf6a665d0fac02ce03e9d3f04f6b46cff38c5f6348ea1caeef1706b807646b803711f55712eed81664309ac826165f70394
6254ac1bead60f90a0edbc9ebb11898b706b807646b80371978a16b13655fe5fa6fcc01e629c6e46706b807646b80371dc0f36563b263c1fe278d2babee8eb06
b2ffa67740ccf7116f1f240f9cc8ca6e706b807646b80371132968115c126500097b19d4c2d9119d706b807646b8037101cbea12ad3dd53b09ac826165f70394
68060a1582a7a49d8a6964f22fb389aa27920222bf9105df2935350fa16e7f91c6696dddf7dbcb67239bdbe658d21d003fa1581d1a600e96bcb8778e5a191662
c5e5d9cd5daf94158b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
*******************************************************************
1e7e75f62a07f7b11a3654f908c2bb013aa2834d09101bc547f3e73fa04e71d0d864ebdf78a436108b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
262b99977648e9d16c5e49ef621538cd706b807646b803715992797124f0124c333cea9549bfb1ed706b807646b80371d209861ab213704e01fc66cb47a60b11
b27e2e819491226c0e8f570a764b71b1b61718b66f0797757ad042da0e82a8d78ba7fe822aeaeae443c740a2312352378b74cc8cf438b7017b9407c104a3fa6d
b2ffa67740ccf7116f1f240f9cc8ca6e706b807646b80371132968115c1265000650ef57a411cfd062d6bdea024861df71a419df3b9cd2e17eb34759a160c424
68060a1582a7a49d6f1f240f9cc8ca6e706b807646b803712935350fa16e7f91097b19d4c2d9119d706b807646b803713fa1581d1a600e96bcb8778e5a191662
c5e5d9cd5daf94158b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
*******************************************************************
d7072740a938f0e737271f6a045506e06194f00f2092c89f7b5b423054b7efee91c26ffb23dc55bd35dee6b9330493134e5235a4865526b9b510bf667672040b
7cafa52502dfe5098b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
b10eccc2ae3b00d8c3872919f6f638ea8c450f0ea0259c5cbdd97c407fe42a54073cd864765286e31a05b145553433318520e268a31fc5ffd7acbf21c6552dd3
e039946fcb76ed7e6fb2315172cc0e50b6721324af5f33cc8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
d7072740a938f0e74a43d4b3f8805fff1ddadd8c1f5214a4275aa0b71223dd186423b436d0b80ef893c50cf5fa8d72419d71b24b6f622a10d3e9d0a2147426cc
*******************************************************************
07673128d177c6cb752e046512a2b14f4f08413eece32388526e666217db2feb1c403045460c978014adac008e277ad86915eb505e8a3b3cfb12c08ee2c37ec0
*******************************************************************
$CDNENCFINISH
.ENDS n36306
*$
**********************************************************************
**********************************************************************
*                                                                    *
*   n36307   -  PSpice Model                                         *
*                                                                    *
*   n36307 is the HS die silicon model for use with 86330q3d         *
*                                                                    *
**********************************************************************
**********************************************************************
* SUBCKT Definition:  1=D  2=G  3=S
**********************************************************************
.SUBCKT n36307  1 2 3
* PARAMETER (local) DEFINITIONS SECTION
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
2cfd781695004e385100148e3d6e300d17b7681b2e59087462d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a96f3b666d9ed3040f
2cfd781695004e387bc7ce494a63b95cab4f8f49c9687b8980fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
2cfd781695004e38126b113ea1f9ad80423ac9b346247ddb60c5ac4de13f4064ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
2cfd781695004e383edbcd936276c8eb36492751f9e6eec919842dc9a1099cd50399937abc26ad30c3444eda896b7868ed857e222a29377b9380942fd2fefa16
2cfd781695004e38444ffe5a14ddde18e488c08cb15a478773bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
****** MODEL SUBCIRCUIT BEGINS HERE     ******************************
1387a7647ddaf4b444ba8c84c92e471c90b8469c307059f0743db0b1d721bf3b93e9a193d756852ef492ccad24701ddac2ec0d54e1fbf00c21ee64457ea555af
13daf902c18c20b08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
d3ae90bb1cd66be0e04afeef43cc7d7162d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
cbe37d5098e0c17824b629fad7d83f95198530b6d3d711d68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
6401eb28bd845c08b1fface195ae7535ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
f569dfd879b57476891e999cbc8ead6639859341766fc92cf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
7a13c2b4abc7a0c32a73071912eabad1ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
1bf2775e5d19f4613cebfa9bcb456bff39859341766fc92cf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
35a1ca33872f2041c6619b7646f07228049104bb5d4ca56dbe401a404cd83ba166fa3ae85270d16309f12bfdd001bf4dc2ec0d54e1fbf00c21ee64457ea555af
13daf902c18c20b08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
3ebc5ddc64c3d282562cd66acf34399062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b324271c0280911f7df87e9386ba9e8f62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
* Note:  gate oxide capacitance included in NMOS below
22118ccc9a4693cbbb823fe98a97c9a6ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
5b8be7694daebfb6b95dbd4ca0a9140ccd0ee77ce9d3a74076617f42cd5d956bf04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
15aa5a803ed33c3095e6484c921cd1d9a722a406594f2665be4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
5cc23a905735a528a38cbb9f2df12ddaf09d6d13bbe7c04dbe4b8e5d291eed266915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbd946b25c2e2c9cf6
*******************************************************************
1e7e75f62a07f7b186e471729bc5541749b5e96410c30f2547f3e73fa04e71d0c24394b0aefd2664706b807646b80371ba80e3b7e443da4b4f85a241c9207b84
262b99977648e9d16c5e49ef621538cd706b807646b80371d3a99143ac7ecc476d570604c7927115f80c4c8e2b766bd8824901d9f53d509df4c83cab6b9aced6
b27e2e819491226c0e8f570a764b71b1b61718b66f0797759c23c515e4041152867b079d0aa545d908e79cbf8de54de39a283b42b20f2dfbd4a932e5ff86e647
809d1592585346e42410f9b01f28bfc2706b807646b80371401e692c311d9e41d1544f4c413476b8706b807646b80371c3be9dd39875721b6b8f064b73f0f573
a284042cd791aa6e58a99dbe66ab556b706b807646b80371ea35a63cd16a7017fe670db4bdff8f92706b807646b803718c2889ca49ca0fe35a9a836056bc521f
3b1feb6bf520a792a25d0694caf72ab8ac8304d24e962dc1bb29955bae8f226fdc4526f415bd9a3fb585b96681e0ca9bfe3ce9cf33d8558c68957789b47fb3f9
4134e00fa366ca83c8d4473d80f8ea33ac8304d24e962dc139b302d18fa67a4258531011761b328da84ecbc7159c51adad084f03a18c1696f62496a6a101fce4
9e13f6a7b30c0d581cd1d6bb2ab26f21706b807646b8037134c64911cb9a3b9ae3568e8b165a35ba706b807646b8037128b2f6472235ee1ed9cd054cffe4113f
ed483728f87a2ff56915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
7b0faa21729cd1dcc65fa3fd5d6e3745706b807646b80371e84c4e9059d274e77a74c1a9b086f5a93421bf8d63a79fc975ae2546e9b9532925bae6d262f7a4f8
5f57011c64ecdeb2e30dea4b4d29e81b706b807646b80371d01a699e884848be787f0235f323548f706b807646b80371c5ed5780386810ae655e130736f46d73
41076da6468fadded813ef29de50e822706b807646b80371e80dcfcbc57bfea854f0b55506f3dab9706b807646b803718b03d7c2720630032e80e42bd2ee1bc1
03dc106fabbcecab6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e7975befcddf1bc8d446e9c238acb2ba0
f8877d765eca4de0592fe1a7ff3cff1a706b807646b803712b20e00307d47b5ee3b5b258cb2aee5c706b807646b80371bb98c84c0bea3b3eb4537737a844a535
1b56e1e057d96a20716a434086c83e8fa665d0fac02ce03e9d3f04f6b46cff383671764b692e1a39706b807646b803711f55712eed81664309ac826165f70394
6254ac1bead60f90a0edbc9ebb11898b706b807646b80371978a16b13655fe5fa6fcc01e629c6e46706b807646b80371dc0f36563b263c1fe278d2babee8eb06
b2ffa67740ccf7116f1f240f9cc8ca6e706b807646b80371132968115c126500097b19d4c2d9119d706b807646b8037101cbea12ad3dd53b09ac826165f70394
68060a1582a7a49d321f85fcffba6c9a27920222bf9105df2935350fa16e7f91c6696dddf7dbcb67239bdbe658d21d003fa1581d1a600e96bcb8778e5a191662
c5e5d9cd5daf94158b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
*******************************************************************
1e7e75f62a07f7b11a3654f908c2bb013aa2834d09101bc547f3e73fa04e71d0d864ebdf78a436108b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
262b99977648e9d16c5e49ef621538cd706b807646b803715992797124f0124cfa594674836cd821706b807646b80371d209861ab213704eece0fa1278d1059f
b27e2e819491226c0e8f570a764b71b1b61718b66f0797757ad042da0e82a8d7871622c33248692eed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
b2ffa67740ccf7116f1f240f9cc8ca6e706b807646b80371132968115c126500097b19d4c2d9119ded857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
68060a1582a7a49d6f1f240f9cc8ca6e706b807646b803712935350fa16e7f91097b19d4c2d9119d706b807646b803713fa1581d1a600e96bcb8778e5a191662
c5e5d9cd5daf94158b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
*******************************************************************
d7072740a938f0e737271f6a045506e01f116e5ac7e8b149378837f1b323cde952ae1caf42661b4d35dee6b9330493134e5235a4865526b9b510bf667672040b
7cafa52502dfe5098b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
0d6f60639959cf60c3872919f6f638ea154202d4ab20f4655fc5f1ba0b28c6660db872e82ffb3e3b1a05b145553433313c09e066d8855370d7acbf21c6552dd3
e039946fcb76ed7e6fb2315172cc0e50b6721324af5f33cc8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
d7072740a938f0e74a43d4b3f8805fff12e6587564d7b4f1275aa0b71223dd186589ec310e2fb4d893c50cf5fa8d72419d71b24b6f622a10d3e9d0a2147426cc
*******************************************************************
07673128d177c6cb752e046512a2b14f4f08413eece32388526e666217db2feb1c403045460c978014adac008e277ad86915eb505e8a3b3cfb12c08ee2c37ec0
*******************************************************************
$CDNENCFINISH
.ENDS n36307


*$


* PSpice Model Editor - Version 16.0.0
*$
.SUBCKT AND2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a911751d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS AND2_BASIC1V
*$
.SUBCKT AND3_BASIC1V A B C Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a91175124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f51d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS AND3_BASIC1V
*$
.SUBCKT AND4_BASIC1V A B C D Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a91175124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bb1d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS AND4_BASIC1V
*$
.SUBCKT NAND2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a91175c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NAND2_BASIC1V
*$
.SUBCKT NAND3_BASIC1V A B C Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a91175124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NAND3_BASIC1V
*$
.SUBCKT NAND4_BASIC1V A B C D Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27aba23a2c92fdb02c4373bf76c56446ed39a9a3702383776c53
ce312808b0a91175124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5124860adb088b20273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bbc4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NAND4_BASIC1V
*$
.SUBCKT OR2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a911751d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS OR2_BASIC1V
*$
.SUBCKT OR3_BASIC1V A B C Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f51d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS OR3_BASIC1V
*$
.SUBCKT OR4_BASIC1V A B C D Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bb1d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS OR4_BASIC1V
*$
.SUBCKT NOR2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a91175c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR2_BASIC1V
*$
.SUBCKT NOR3_BASIC1V A B C Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR3_BASIC1V
*$
.SUBCKT NOR4_BASIC1V A B C D Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab989d941548be479d73bf76c56446ed39a9a3702383776c53
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bbc4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR4_BASIC1V
*$
.SUBCKT NOR5_BASIC1V A B C D E Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161ef0070e980448d49ce5ec34e6f8ad1ca4f07b1c061ae9cfeab0e2d7cadb195efd4198695988ed1bb8b74cc8cf438b7017b9407c104a3fa6d
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bbe22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
bdac9a78f852a4f3c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR5_BASIC1V
*$
.SUBCKT NOR6_BASIC1V A B C D E F Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161ef0070e980448d49ce5ec34e6f8ad1ca4f07b1c061ae9cfeab0e2d7cadb195efd4198695988ed1bb8b74cc8cf438b7017b9407c104a3fa6d
ce312808b0a91175e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
49482642e74b34f5e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
558aa0970ce534bbe22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
bdac9a78f852a4f3e22c09012d03f80973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
6a60a2b3c07c62b9c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR6_BASIC1V
*$
.SUBCKT INV_BASIC1V A  Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab1e9e9577d905ee24ddf7ad811d6a72c444eb3bb0fc4b8a93
9ee3082acb32f34aed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS INV_BASIC1V
*$
.SUBCKT XOR2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161492f206f537e28b38492e52ca99071372a4b8dedaaff0e2c27bb8ad2fa403e2b164ffd829dfc9575ddf7ad811d6a72c444eb3bb0fc4b8a93
ce312808b0a911751d30254c6c3ade365741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS XOR2_BASIC1V
*$
.SUBCKT XNOR2_BASIC1V A B Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161492f206f537e28b38492e52ca99071372a4b8dedaaff0e2c27bb8ad2fa403e2b164ffd829dfc9575ddf7ad811d6a72c444eb3bb0fc4b8a93
ce312808b0a91175c4475f08bdea21f15741e5db7e96aaea8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS XNOR2_BASIC1V
*$
.SUBCKT MUX2_BASIC1V A B S Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161492f206f537e28b38492e52ca99071378fef95ad867776d986d7aaf828690538bf1ee911780421dd6915eb505e8a3b3cfb12c08ee2c37ec0
d5c1d990d4a5ccdb03d5eef6b3061dfa73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS MUX2_BASIC1V
*$
.SUBCKT INV_DELAY_BASIC1V A  Y PARAMS: DELAY = 10n
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161b7a8d0a5fa27600f87c337a6226f9c259ce2376dcef929e055e2d3dce1717d719697193234a3017f73bf76c56446ed39a9a3702383776c53
933bd4b4ee0a4eaeed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
bd9831b9881f0b92004c220067cfdabf57e2c5aa808513706915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99cb3fa3ad4040ee39d350e60ca2338a43558a6d1f49bc89ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
f305b7cfa0765161c36180965553170d8da13727b91264449ce2376dcef929e07d4a1829490ab8db27bb8ad2fa403e2b040397452ddd04155a97c8100a7f5192
9ee3082acb32f34aed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
8d3568177ac8ace9a0338d780f826fc662d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
042d1e8ae349b80f5801d29f353ff668ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f62c8b4f8e886a69cc
$CDNENCFINISH
.ENDS INV_DELAY_BASIC1V
*$
.SUBCKT BUF_DELAY_BASIC1V A  Y PARAMS: DELAY = 10n
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa0765161b7a8d0a5fa27600f87c337a6226f9c259ce2376dcef929e055e2d3dce1717d719697193234a3017f73bf76c56446ed39a9a3702383776c53
933bd4b4ee0a4eaeed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
bd9831b9881f0b92004c220067cfdabf57e2c5aa808513706915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99cb3fa3ad4040ee39d350e60ca2338a43558a6d1f49bc89ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
f305b7cfa0765161c36180965553170d8da13727b91264449ce2376dcef929e07d4a1829490ab8db27bb8ad2fa403e2b040397452ddd04155a97c8100a7f5192
933bd4b4ee0a4eaeed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
8d3568177ac8ace9a0338d780f826fc662d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
042d1e8ae349b80f5801d29f353ff668ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1fa3e5af8a9f0d59f62c8b4f8e886a69cc
$CDNENCFINISH
.ENDS BUF_DELAY_BASIC1V
*$
.SUBCKT BUF_BASIC1V A  Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751893d7ec53d9f27ab1e9e9577d905ee24ddf7ad811d6a72c444eb3bb0fc4b8a93
933bd4b4ee0a4eaeed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS BUF_BASIC1V
*$
**Set has higher priority in this latch
.SUBCKT SRLATCHSHP_BASIC1V S R Q QB
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc249a0b346cfeb7a8aee7af706d286b8b361830ae1f2a413b17a9af17d7769a2bcdfd7acbf21c6552dd3
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b39212aa4361a7de9e97ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de1adbce7254a8ccba480fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa767080305345996932e974031f2ece18280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08ef8e5128bbe27bfd2c
8f7b8724f31a9e8c1250a7e9a95e2aa381ed1a17eaffcba773bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS SRLATCHSHP_BASIC1V
*$
**Reset has higher priority in this latch
.SUBCKT SRLATCHRHP_BASIC1V S R Q QB
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24918f1e062ef55a242af1b6d78a26c00872c2a5798878066b49af17d7769a2bcdfd7acbf21c6552dd3
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b39212aa4361a7de9e97ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de1adbce7254a8ccba480fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa7b47141f0f87379b062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
8f7b8724f31a9e8c9bb209fe8097ada262d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
cb3de6a18d5d6014341eeb2a089c5b4f80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS SRLATCHRHP_BASIC1V
*$
**Reset has higher priority in this latch and active low set and reset - basically NAND based SR latch
.SUBCKT SBRBLATCHRHP_BASIC1V SB RB Q QB
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24909bbe8dd12e94074cfdf74b4198081a0ff507e01fe1ffea7cb09da6dde53e4e5ed39ea6b8106f78c
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b39212aa4361a7de9e97ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de1adbce7254a8ccba480fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS SBRBLATCHRHP_BASIC1V
*$
**Reset has higher priority in this latch and active low set and reset - basically NAND based SR latch
.SUBCKT SBRBLATCHSHP_BASIC1V SB RB Q QB
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24956921f5b7804ee684e4a831e2a781a75d75465cefb0b0b029b7057a214a14dbfed39ea6b8106f78c
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b39212aa4361a7de9e97ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de1adbce7254a8ccba480fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS SBRBLATCHSHP_BASIC1V
*$
.SUBCKT DFFSBRB_SHPBASIC1V Q QB CLK D RB SB
***Set has higher priority in this
** Changed the delay from 7n/10n to 15n/20n to help larger time step simulations
**Faster flip-flops require a a smaller time step to simulate
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
e347113957ea6865794f28b54474bef138d847730d715c66a48f4886f5e648f71933952b4dcad44c7980309da51cc49d59d51a6aaa99d5782bb0da26e91d20fe
1e3cbcba78a2571717c616a6bb942482b8e5f1c1d9b7fc962d3711465512234c1b58fcc31687397c6915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24956921f5b7804ee684e4a831e2a781a7577955cbe1d3455d964d27582d4f28f719a4b29c3b5d68e76
624fde9c288b3ae2644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
c2b7a0b474b4bcc083b19b9f68334754dbb6b6ac355aa998e71f71e187584171f04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b3929c99a6f8ecce3483903bfb975c9062585441d228f64798f82fdbf39023f863b5e5d5c6a1b5a1b63a5a97c8100a7f5192
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de197607e8fde09e5ae80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa7c9380a751924b9b2ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
8f7b8724f31a9e8cbe63f4e3bfd183b0644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS DFFSBRB_SHPBASIC1V
*$
.SUBCKT DFFSR_SHPBASIC1V Q QB CLK D R S
***Set has higher priority in this
** Changed the delay from 7n/10n to 15n/20n to help larger time step simulations
**Faster flip-flops require a a smaller time step to simulate
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
e347113957ea6865794f28b54474bef138d847730d715c66a48f4886f5e648f71933952b4dcad44c7980309da51cc49d59d51a6aaa99d5782bb0da26e91d20fe
1e3cbcba78a2571717c616a6bb942482b8e5f1c1d9b7fc962d3711465512234c1b58fcc31687397c6915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc249a0b346cfeb7a8aee7af706d286b8b36118f1e062ef55a24264d27582d4f28f719a4b29c3b5d68e76
624fde9c288b3ae2644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
c2b7a0b474b4bcc083b19b9f68334754dbb6b6ac355aa998e71f71e187584171f04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b3929c99a6f8ecce3483903bfb975c9062585441d228f64798f82fdbf39023f863b5e5d5c6a1b5a1b63a5a97c8100a7f5192
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de197607e8fde09e5ae80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa7c9380a751924b9b2ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
8f7b8724f31a9e8cbe63f4e3bfd183b0644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS DFFSR_SHPBASIC1V
*$
.SUBCKT DFFSBRB_RHPBASIC1V Q QB CLK D RB SB
***Set has higher priority in this
** Changed the delay from 7n/10n to 15n/20n to help larger time step simulations
**Faster flip-flops require a a smaller time step to simulate
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
e347113957ea6865794f28b54474bef138d847730d715c66a48f4886f5e648f71933952b4dcad44c7980309da51cc49d59d51a6aaa99d5782bb0da26e91d20fe
1e3cbcba78a2571717c616a6bb942482b8e5f1c1d9b7fc962d3711465512234c1b58fcc31687397c6915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24909bbe8dd12e94074cfdf74b4198081a02f2603dd7679f7f20c965cdf587c9d6f9a4b29c3b5d68e76
624fde9c288b3ae2644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
c2b7a0b474b4bcc083b19b9f68334754dbb6b6ac355aa998e71f71e187584171f04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b3929c99a6f8ecce3483903bfb975c9062585441d228f64798f82fdbf39023f863b5e5d5c6a1b5a1b63a5a97c8100a7f5192
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de197607e8fde09e5ae80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa7c9380a751924b9b2ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
8f7b8724f31a9e8cbe63f4e3bfd183b0644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS DFFSBRB_RHPBASIC1V
*$
.SUBCKT DFFSR_RHPBASIC1V Q QB CLK D R S
***Set has higher priority in this
** Changed the delay from 7n/10n to 15n/20n to help larger time step simulations
**Faster flip-flops require a a smaller time step to simulate
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
e347113957ea6865794f28b54474bef138d847730d715c66a48f4886f5e648f71933952b4dcad44c7980309da51cc49d59d51a6aaa99d5782bb0da26e91d20fe
1e3cbcba78a2571717c616a6bb942482b8e5f1c1d9b7fc962d3711465512234c1b58fcc31687397c6915eb505e8a3b3c33ef52353febd1f220ba217fa27494f5
08e147163f37b483eb1553db51121b0af03ffeaf6f4cc24918f1e062ef55a242af1b6d78a26c00879055549affe647300c965cdf587c9d6f9a4b29c3b5d68e76
624fde9c288b3ae2644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
c2b7a0b474b4bcc083b19b9f68334754dbb6b6ac355aa998e71f71e187584171f04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
a405048fcac30c1a338602ff93fff92d62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
b75a50bb44e3b503f2667b5cb330c5cf12000876fc7937f7ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe32fb8e6d82984fc1f68b06386d7b2f79a
1033be605ac86fd802147ff4d5c4cb2f895d090a759f83318b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
4d7ee7dde33e93874d2f23a30635e4366915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
7b341edfa7445b08bd6fc2e97e23189d303d7240d8c3139d6915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
99fafaa2580fb990086c1f20d6d180eb36806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
b8c0b98b8ee14d0e86fb6fea0644b3929c99a6f8ecce3483903bfb975c9062585441d228f64798f82fdbf39023f863b5e5d5c6a1b5a1b63a5a97c8100a7f5192
7e2980978c86958c3c22444f975fafc280fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
161224ee3eeadb9c8492e52ca99071370aa8feaa9dcff151057d265e60bc684b84d9bb7728971e45ed857e222a29377b14aee5f82b16b767a53ed4fb58cd5d2b
04db544825bf7de197607e8fde09e5ae80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
97c9333151ea8fa7c9380a751924b9b2ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
8f7b8724f31a9e8cbe63f4e3bfd183b0644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
cb3de6a18d5d601472130360ca424be562d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
d7072740a938f0e76796778f313a81b5bcf1ee82bdd45fd86d0ad17b3ef49a3d2ed4e03f3e56f24b32b39d3050b302d280fa21721bf3358cc4169e4a88b5de56
$CDNENCFINISH
.ENDS DFFSR_RHPBASIC1V
*$
.SUBCKT DFFSBRB_RHPBASIC1VVxxx2 Q QB CLK D RB SB
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
0396f539ca92147d57a2d954b5055c78ff5b4ecc92f3c4136ba07ab578b94b9315e672de8a85df84fde82b3677c6a11ec11c2062aece1f332286150040758a84
a978e94c36773adb4ac7590e81b8b7fe282c6e10dcffb68c85c227248672f89b50f00e03b07d40457e72cfc55f390f1f3adb303f5db25bc503b0837954bde256
22d19f90c399e00ded857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
2945e767cc1052a3c058a76726120dbf71f52ef20542de6443706c6781e88dd56836447af54d14090c994f1d777bc8e5ed857e222a29377b9380942fd2fefa16
a978e94c36773adb4ac7590e81b8b7fe282c6e10dcffb68c85c227248672f89b0b663d2bae9992e97e72cfc55f390f1f80472ae340292c1103b0837954bde256
22d19f90c399e00ded857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a022c9b4089f2aa3283508d19ff419fb587f
bb80ebdc847f079a63717d323a8bd56aa48f4886f5e648f7ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
3637782305084aad5e58a4711fa34dc1dc4d3e8d456b5b64b91f6756c247f62c8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398f317f2de0bd9ffbe
538cf038f20f7f797961a41b1a118afaa48f4886f5e648f7ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
6cc754a414c3ec967961a41b1a118afaa48f4886f5e648f7ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
0de082d7aaf8348a5baf4eb20ab697209ab22aaa94d8499e2191821dd460f2248bfd91f88313a65962d6bdea024861df71a419df3b9cd2e17eb34759a160c424
$CDNENCFINISH
.ENDS DFFSBRB_RHPBASIC1VVxxx2
*$
.SUBCKT DLATCHSR_PS1 D CLK Q0 QN SB RB
+  PARAMS: vhi=1 vlo=0 vthresh=0.5 tplh=1e-9 tphl=1e-9 tr=1e-9 tf=1e-9
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
abddc8f1b1c320096044af6e2c9f213b1cf484586c5b834452c47937a970f2d74806f38dfed245548b74cc8cf438b701ea09ec4bf584f8dd55869a830df61378
a978e94c36773adb4ac7590e81b8b7fe282c6e10dcffb68c85c227248672f89be5d1361524860fbded3fe434838c12cfdb927fe7f2ae9c00800a01cc1bdb843c
9b65bac9ecb5f6aec1e35104f25f8b0073bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
ff644bacb164bd15964067500402814c6baa4c351fc5e3adcb9b72e106d1d63573bf76c56446ed39c27a29c2d535fd4ea444f95e85eea42155a6f3f1d348a0ee
7c964f6453abbae954588f17103cc829a74fe0b4f4ce2af9a48f4886f5e648f7ed857e222a29377b14aee5f82b16b7673d4db86b42817e2bf411d12d7ec6c2f4
c94eb5aabc7a5cfe64146fdf1779d397fa460eccc75cda6deb1f486074fe0c28ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
3690e7acd67ee7d33511aefda81833ee726d9a7f6b37359cb27cc86ab8fb764a80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd5469306ad371de54
cba19b3e6911e6dac68dcb01828c2c574ac5ddcf254124727662f9e929a451eeb27cc86ab8fb764a80fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
16d01f52c0c1b16ae504ac4df1b1e2bc9733fa0a03265685a873c24146caa13062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
b23966fe8e7921c4988ba3fc13166d49d8286d136f179c49a873c24146caa13062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
a19132db4faf0e2553aadc974be762875bf56a7c0e781c9d6f3096029d06b975a5dd93e2580e537f73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
5b52b71f43a037c6fd70c76153b2d299a5dd93e2580e537f73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
***X9 Sint1 Setlogic Sint OR2_BASIC1V
****X10  Rint1 Resetlogic Rint OR2_BASIC1V
$CDNENCFINISH
.ENDS DLATCHSR_PS1
*$
.SUBCKT DLATCHSR_PS2 D CLK Q0 QN SB RB
+ PARAMS: vhi=1 vlo=0 vthresh=0.5 tplh=1e-9 tphl=1e-9 tr=1e-9 tf=1e-9
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
abddc8f1b1c320096044af6e2c9f213b1cf484586c5b834452c47937a970f2d7bd70f954bb2c8c96ddf7ad811d6a72c40790ffaf43e25844c4d2097fcab0f49a
a978e94c36773adb4ac7590e81b8b7fe282c6e10dcffb68c85c227248672f89be5d1361524860fbded3fe434838c12cfdb927fe7f2ae9c00800a01cc1bdb843c
9b65bac9ecb5f6aec1e35104f25f8b0073bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
ff644bacb164bd15964067500402814c6baa4c351fc5e3adcb9b72e106d1d63573bf76c56446ed39c27a29c2d535fd4ea444f95e85eea42155a6f3f1d348a0ee
7c964f6453abbae954588f17103cc829a74fe0b4f4ce2af9a48f4886f5e648f7ed857e222a29377b14aee5f82b16b7673d4db86b42817e2bf411d12d7ec6c2f4
c94eb5aabc7a5cfe64146fdf1779d397fa460eccc75cda6deb1f486074fe0c28ddf7ad811d6a72c40790ffaf43e25844402a22a00a175fe31c80df6ba8cb4d47
3690e7acd67ee7d33511aefda81833ee726d9a7f6b37359cb27cc86ab8fb764a80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd5469306ad371de54
cba19b3e6911e6dac68dcb01828c2c574ac5ddcf254124727662f9e929a451eeb27cc86ab8fb764a80fa21721bf3358ca6de71685bf58c903a5dc079a48bd340
16d01f52c0c1b16ae504ac4df1b1e2bc9733fa0a03265685a873c24146caa13062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
b23966fe8e7921c4988ba3fc13166d49d8286d136f179c49a873c24146caa13062d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a615ba3ed11d2389294
a19132db4faf0e2553aadc974be762875bf56a7c0e781c9d6f3096029d06b975a5dd93e2580e537f73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
5b52b71f43a037c6fd70c76153b2d299a5dd93e2580e537f73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
***X9 Sint1 Setlogic Sint OR2_BASIC1V
****X10  Rint1 Resetlogic Rint OR2_BASIC1V
$CDNENCFINISH
.ENDS DLATCHSR_PS2
*$
.SUBCKT NORLATCHDFF_PS SET RESET Q0 QN PARAMS: vhi=1 vlo=0 vthresh=0.5 tplh=1e-9 tphl=1e-9 tr=1e-9 tf=1e-9
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
1f32d041af08515ad7070c5fa5f708f81e6056a43023a69462d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a96f3b666d9ed3040f
16a6899257d114c6d7070c5fa5f708f8e26b1054de4177ca62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a96f3b666d9ed3040f
c3dd5b5fc815d5491cc283117763bd2732273240e56ef04c55cc7113ef7d91bdc25420ed8957389351045afd8f3f23982414ad3f96a2b449017b011f6d57fcfa
024c16587eeb9d355ed675620634412b180865aa314321c1d5e0deeab85ec3dc77387bc0bba0a96e73bf76c56446ed39c27a29c2d535fd4e755b4380fba48b25
25a93b8a68c28939b8f058f964dbea42266bfb5b138f20b19456dd01a5954e548743172692865944b573d8e00b32e08ebb4d5d880284260c91301b0d831affca
bc557f4f0b62c9a9b4428d603bd51a53f033cbe1442b49a9b976213f12230533aa0ec03329b1d41433778b5e19c8d4e3c612182fe29e690d5a97c8100a7f5192
733c41074305b5a95b9f97e31a6d9c8612aa4361a7de9e97644126c9831a96bdf04163af94c95a1d0d3a4073c77cf923dc361e602ca60976ef88b43b2e5ecd8a
bba3d5a11127e656dde6c88d33167b8112aa4361a7de9e97ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
$CDNENCFINISH
.ENDS NORLATCHDFF_PS
*$
.SUBCKT NOR2_PS Y A B PARAMS: vhi=1 vlo=0 vthresh=500e-3 tplh=1e-9 tphl=1e-9 tr=1e-9 tf=1e-9
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
b1e1a75a4c03144fb84942cebd8cf2b68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
383821663e4954c2f610485492ce8d1980fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
6b5d5a08a2b08391b84942cebd8cf2b68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
ca3c8af328efcba6f610485492ce8d1980fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
f0a3943a524b95e16bcb608151f4536673bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
5843b7df5950ebb53bfc9ee8dc6e0fd25414ce0c3c28bd7fd1150c70c992e76f2395ba5dcc96121f32cf6bdf8be6e9e830d880300d5bb3510c8cfd52bfe4b3c7
4bbf5fa8614861d08b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f8070ecac8716a4aa4ae489193d39b540
1830c2657ad72cfd80caf75d9556d4e836806a8e381bf9a0f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b86110972015b4a108
e683a3d374597388319394d2970bb1aebf0e8aeac1ee4acf1933952b4dcad44c4d985589162d35b85192a1f4ea15cca8c6314e3c21f3975457088b21e284207f
59696ce43217c78a489d02fabd515895ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
50ff5937e1f4aec7088a4decac19c24efa15b6f6532689ccbff077c5371b976ad899b67b1514e77c247ce4099c7069888ed9989b4fdbe89c84a603f467791872
b6740db0d75566c15bd9ba46c107a781ee296b5d6cfe99f68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584bc723f2834d23f68
e65068a5529a5a08bc8abe03198c62e2ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
4c1a4bf8a33698824a3bc44e792baa17979added4bba322b45555c45879de233c3b775f7138ddffa8ee54616d1c590f4ddf7ad811d6a72c444eb3bb0fc4b8a93
4acc2604cc13e40087d03543a42c123a62d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
f5ece99b8dc1e922134ba678c3a552ab9286534c194f5bf760129872902b40542852f737f3e1fdd297efe455f1ba5b5566c5e322d06d2953a2713860206d5dfb
5bd9ba46c107a781ee296b5d6cfe99f68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
230c8a132db19d25c306c8e91cade4aa18018bad8db9c9d30c4f3a1c4714b0fa69413a540c7bb72fc3c82ada44c780f2c6314e3c21f397544afce059d1020bbe
e0dfb329be65daf28f98c50ec84605b673bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
bd6fe760313481fff7307a8bcc75d233ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
d1579de13894cc532e865137b41094437d1b42c81d7f147d8795a8d338813804060e5e0af582bfca237b8d7a10235eade71f71e187584171cad25bf5db12395b
f9da05a8e6a65298826d20fdd211253fed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbc002d19ceb77a0227332f86ebd489748
d78f19d4db97b9b7b84942cebd8cf2b68b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS NOR2_PS
*$
.SUBCKT PSW_PS D G S PARAMS: RONval=10k VTHval=0.7 VCHARval=0.01 CGval=0.01pF CDval=0.01pF
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
3f510a0fa0d9a58d00037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
4fee993ae8eff14300037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
c8baedcc8773edc600037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
36e77ffbd2e958de9ce28abedde281fd73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
4c3141c46a36e1abda49105010470d0173bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
bcc2b5d8d2a44ed3e36ada7603e37bde979added4bba322b584a1251b11bb09b8577b07d1241b40e26d29dc8994456ec13ba82e50acd77deee626c3c1261d425
5a8ca3732b7d40643f730f3e2357fdcd72cc4e0395929afecaa5e0711288816a3e3bed9e00fb4633714f855d3587b318000fc12d735d5beb69ba81bc9f61e2f4
ceaf4f6c775c0b0150a36120f822a26cc28bd7eced7ae73273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
$CDNENCFINISH
.ENDS PSW_PS
*$
.SUBCKT NSW_PS D G S PARAMS: RONval=10k VTHval=0.7 VCHARval=0.01 CGval=0.01pF CDval=0.01pF CSval=0.01pf
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
3f510a0fa0d9a58d00037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
4fee993ae8eff14300037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
c8baedcc8773edc600037464c659791973bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
36e77ffbd2e958de9ce28abedde281fd73bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
4c3141c46a36e1abda49105010470d0173bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
8f1407e2c16ee8e828717dfc8175393473bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920736773acebe3f8d53d23d74009f155f7
***EEXP F1 0 VALUE={LIMIT(((V(G,S)-VTHval)/VCHARval),-80,80)}
bcc2b5d8d2a44ed3e36ada7603e37bde979added4bba322b7236a99fbbbba11e632a2f36d939f491632a2f36d939f491f12736b1ad219720ee626c3c1261d425
6344dda27888449d3f730f3e2357fdcdd88055922e5b0740caa5e0711288816a3e3bed9e00fb4633714f855d3587b318000fc12d735d5beb69ba81bc9f61e2f4
ceaf4f6c775c0b0150a36120f822a26cc28bd7eced7ae73273bf76c56446ed39c27a29c2d535fd4ea444f95e85eea421e624fc2223ab3920f0189eec88ecdc90
$CDNENCFINISH
.ENDS NSW_PS
*$






*$
.SUBCKT COMP_BASIC1V INP INM Y
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
324d0b28bd3976fec3fa3d1e401a4503c7cd3c6de157579e2a235350161d1bcb644126c9831a96bdf04163af94c95a1d0d3a4073c77cf9236dc1cba06b961a0c
31a245cc4f39b9f137f223f6cbbe63d162d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
3b7f5ebe940d64624170694978eb4cf88b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
b076ff8d9576189163285b2908224391f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
$CDNENCFINISH
.ENDS COMP_BASIC1V
*$
.SUBCKT COMPHYS_BASIC1V INP INM HYS OUT
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
9132b7121104d4358be44c41ab888f41b6e3a1568843d867ed857e222a29377b14aee5f82b16b7673d4db86b42817e2b94029deb845b63dbfa609432f74b4cf3
70d49a25931fcad5af5f0f227a33dfc56b574213c15e8d89a3a038b03e03563d54d03668c743d1a6bb77e20fe987edd8ed857e222a29377b9380942fd2fefa16
d1579de13894cc53749d13634498f34b2814ec203481f38f6485690991963efc688dc2cfc32ec3a971a7af633826d31662d6bdea024861df2dd112e4aa362c02
c985c90e830fff9457e2c5aa808513706915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
1fdb31c906bbcd7763285b2908224391f04163af94c95a1d0d3a4073c77cf923dc361e602ca609762950f096084b66b860df248993afc75fcc58c2ffb82de3eb
13142c038a62aa150aa66cfdd7abddd762d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
$CDNENCFINISH
.ENDS COMPHYS_BASIC1V
*$


*$
.SUBCKT LDCR 1 2 PARAMS: L=1u DCR=20m
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
3ef58a3cc4ced0ee35574dcb5fb4fe8080fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
48d1201f22a6f79d5d9f033cb3c2bb5462d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
$CDNENCFINISH
.ENDS LDCR
*$
.SUBCKT CESR 1 2 PARAMS: C=10u ESR=2m ESL=1n
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
3cea00e3e3d5df881915be8fc72309be80fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
48d1201f22a6f79d0d80c60f3da72cbc0b84675c82dbaa586915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d4812c93bd6c982cd5
8450d0214889964a118d53f5ccda89c962d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b5872426f8a8ef40a28
$CDNENCFINISH
.ENDS CESR
*$
*$
.SUBCKT AND2_BASIC_GEN A B Y PARAMS: VDD=1 VSS=0 VTHRESH=0.5
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
f305b7cfa07651615a9037c8c42a602b94aebb18efc1b73c4a0534bc16c6b751d67091752c09698a1541fe9d381cc675621f57e8bf9b586eee626c3c1261d425
ce312808b0a91175dcf306adebf133c01a6c7500361cb5a45652e10015a645e7e71f71e187584171f04163af94c95a1d0d3a4073c77cf9236dc1cba06b961a0c
bd9831b9881f0b92e8f02e93fcf213a880fa21721bf3358ca6de71685bf58c900983ad7c94dcefbd14f1317035ef08efdd67fe27271281584e4e63a74e7b29eb
02f2959404528fbd9ad2dc2e0af5de0e8b74cc8cf438b701ea09ec4bf584f8dd281b4bcb2fc65398d456790f533c7584c8e64aca10a7361f123a3133a745b941
$CDNENCFINISH
.ENDS AND2_BASIC_GEN
*$







.MODEL DD1 D
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
c6d73252edd0ce7a47ebccea066b33f8a262f2beadd5de8083a9e4a7c156932ea67a7ba872982cbd14aee5f82b16b7673d4db86b42817e2bf411d12d7ec6c2f4


$CDNENCFINISH



.model dd d
$CDNENCSTART
eee8c5c7a2bc4b01f045f303678664e7916da0bae22e8cb0bba041dd67c69ce448ea70148a9ac1670c8926c1ac5057c8ccfcd77bf87ca9dc5a97c8100a7f5192
017be2304022735962d6bdea024861df71a419df3b9cd2e10f73aa04b9c40a61ee80317e3f8c42a92e2a580c88a20b581739c5c1ab2d23f214b807900fe3ac5c
39c84b0c9f72e00767286f562e81c2a26915eb505e8a3b3c33ef52353febd1f2ca9826ced64f37cbf69d44061c3450d426dc457f7871e36e5c9ba9c17300437f
*.MODEL D_D1 D( IS=1e-15 TT=10p Rs=0.05 N=.1 )

$CDNENCFINISH
