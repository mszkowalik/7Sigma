.SUBCKT MCP6V11 1 2 3 4 5
*               | | | | |
*               | | | | Output
*               | | | Negative Supply
*               | | Positive Supply
*               | Inverting Input
*               Non-inverting Input
*
********************************************************************************
* Software License Agreement                                                   *
*                                                                              *
* The software supplied herewith by Microchip Technology Incorporated (the     *
* 'Company') is intended and supplied to you, the Company's customer, for use  *
* soley and exclusively on Microchip products.                                 *
*                                                                              *
* The software is owned by the Company and/or its supplier, and is protected   *
* under applicable copyright laws. All rights are reserved. Any use in         *
* violation of the foregoing restrictions may subject the user to criminal     *
* sanctions under applicable laws, as well as to civil liability for the       *
* breach of the terms and conditions of this license.                          *
*                                                                              *
* THIS SOFTWARE IS PROVIDED IN AN 'AS IS' CONDITION. NO WARRANTIES, WHETHER    *
* EXPRESS, IMPLIED OR STATUTORY, INCLUDING, BUT NOT LIMITED TO, IMPLIED        *
* WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE APPLY TO  *
* THIS SOFTWARE. THE COMPANY SHALL NOT, IN ANY CIRCUMSTANCES, BE LIABLE FOR    *
* SPECIAL, INCIDENTAL OR CONSEQUENTIAL DAMAGES, FOR ANY REASON WHATSOEVER.     *
********************************************************************************
*
* The following op-amps are covered by this model:
*      MCP6V11, MCP6V11U
*
*
* Revision History:
*      REV A: 17-MAY-12, Created model
*      REV B: 09-Jul-12, Added MCP6V11U
*
*
*
*
* Recommendations:
*      Use PSPICE (or SPICE 2G6; other simulators may require translation)
*      For a quick, effective design, use a combination of: data sheet
*            specs, bench testing, and simulations with this macromodel
*      For high impedance circuits, set GMIN=100F in the .OPTIONS statement
*
* Supported:
*      Typical performance for temperature range (-40 to 125) degrees Celsius
*      DC, AC, Transient, and Noise analyses.
*      Most specs, including: offsets, DC PSRR, DC CMRR, input impedance,
*            open loop gain, voltage ranges, supply current, ... , etc.
*      Temperature effects for Ibias, Iquiescent, Iout short circuit
*            current, Vsat on both rails, Slew Rate vs. Temp and P.S.
*
* Not Supported:
*      Some Variation in specs vs. Power Supply Voltage
*      Vos distribution, Ib distribution for Monte Carlo
*      Distortion (detailed non-linear behavior)
*      Some Temperature analysis
*      Process variation
*      Behavior outside normal operating region
*
* Known Discrepancies in Model vs. Datasheet:
*      Only analog functions modelled.  CS ignored.
*      Saturation recovery model does not accurately predict recovery time.
*
*
* Input Stage
V10  3 10 -210M
R10 10 11 69.0K
R11 10 12 69.0K
G10 10 11 10 11 1.44M
G11 10 12 10 12 1.44M
C11 11 12 76.8P
C12  1  0 6.00P
E12 71 14 POLY(6) 20 0 21 0 22 0 23 0 26 0 27 0   700N 12.3 12.3 12.3 12.3 1 1
G12 1 0 62 0 1m
G13 1 2 63 0 1u
M12 11 14 15 15 NMI
M14 12 2 15 15 NMI
G14 2 0 62 0 1m
C14  2  0 6.00P
I15 15 4 500U
V16 16 4 10.0M
GD16 16 1 TABLE {V(16,1)} ((-100,-100E-15)(0,0)(1m,1u)(2m,1m))
V13 3 13 -10.0M
GD13 2 13 TABLE {V(2,13)} ((-100,-100E-15)(0,0)(1m,1u)(2m,1m))
R71  1  0 10.0E12
R72  2  0 10.0E12
R73  1  2 10.0E12
*C13  1  2 3.00P
*
* Noise, PSRR, and CMRR
I20 21 20 423U
D20 20  0 DN1
D21  0 21 DN1
I22 22 23 1N
R22 22 0  1k
R23  0 23 1k
G26  0 26 POLY(2) 3 0 4 0   0.00 -177U -177U
R26 26  0 1
G27  0 27 POLY(2) 1 0 2 0  -1.73U 100N 100N
R27 27  0 1
*
* Open Loop Gain, Slew Rate
G30  0 30 12 11 1
R30 30  0 1.00K
G31 0 31 3 4 5.83
I31 0 31 DC 29.5
R31 31  0 1 TC=3.05M,-14.5U
GD31 30 0 TABLE {V(30,31)} ((-100,-1n)(0,0)(1m,0.1)(2m,2))
G32 32 0 3 4 12.5
I32 32 0 DC 31.9
R32 32  0 1 TC=2.46M,-16.5U
GD32 0 30 TABLE {V(30,32)} ((-2m,2)(-1m,0.1)(0,0)(100,-1n))
G33  0 33 30 0 1m
R33  33 0 1K
G34  0 34 33 0 1.77
R34  34 0 1K
C34  34 0 2.83M
G37  0 37 34 0 1m
R37  37 0 1K
C37  37 0 159P
G38  0 38 37 0 1m
R38  39 0 1K
L38  38 39 318U
E38  35 0 38 0 1
G35 33 0 TABLE {V(35,3)} ((-1,-1n)(0,0)(50.0,1n))(55.0,1))
G36 33 0 TABLE {V(35,4)} ((-55.0,-1)((-50.0,-1n)(0,0)(1,1n))
*
* Output Stage
R80 50 0 100MEG
G50 0 50 57 96 2
R58 57  96 0.50
R57 57  0 100
C58  5  0 2.00P
G57  0 57 POLY(3) 3 0 4 0 35 0 0 3.75M 5.00M 10.0M
GD55 55 57 TABLE {V(55,57)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
GD56 57 56 TABLE {V(57,56)} ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
E55 55  0 POLY(2) 3 0 51 0 -800U 1 -56.0M
E56 56  0 POLY(2) 4 0 52 0 566U 1 -45.7M
R51 51 0 1k
R52 52 0 1k
GD51 50 51 TABLE {V(50,51)} ((-10,-1n)(0,0)(1m,1m)(2m,1))
GD52 50 52 TABLE {V(50,52)}  ((-2m,-1)(-1m,-1m)(0,0)(10,1n))
G53  3  0 POLY(1) 51 0  -500U 1M
G54  0  4 POLY(1) 52 0  -500U -1M
*
* Current Limit
G99 96 5 99 0 1
R98 0 98 1 TC=-7.61M,25.6U
G97 0 98 TABLE { V(96,5) } ((-11.0,-8.00M)(-1.00M,-7.92M)(0,0)(1.00M,7.92M)(11.0,8.00M))
*E97 99 0 VALUE { V(98)* LIMIT(((V(3)-V(4))*375M + 62.5M),0.05,1E6)}
E97 99 0 VALUE { V(98)* LIMIT(((V(3)-V(4))*375M + 62.5M),0.00,1E6) *
+ LIMIT(((V(3)-V(4))*400M + 0.00),0,1)}
D98 4 5 DESD
D99 5 3 DESD
*
* Temperature / Voltage Sensitive IQuiscent
R61 0 61 1 TC=2.70M,-7.11U
G61 3 4 61 0 1
G60 0 61 TABLE {V(3, 4)}
+ ((0,0)(500M,61.0N)(1.5,5.6U)(2.5,5.8U)
+ (3.5,6.00U)(4.5,6.1U)(5.5,6.2U))
*
* Temperature Sensitive offset voltage
I73 0 70 DC 1uA
R74 0 70 1 TC=50.0M
E75 1 71 70 0 1
*
* Temp Sensistive IBias
*I62 0 62 DC 1uA
I62 0 62 DC 1000uA
R62 0 62 REXP  49.57961U
*
* Temp Sensistive Offset IBias
I63 0 63 DC 1uA
R63 0 63 25.0 TC=56.1M,597U
*
* Models
.MODEL NMI NMOS(L=2.00U W=42.0U KP=200U LEVEL=1 )
.MODEL DESD  D   N=1 IS=1.00E-15
.MODEL DN1 D   IS=1P KF=14.6E-18 AF=1
.MODEL REXP  RES TCE= 4.20742
.ENDS MCP6V11

