* Resistor
.subckt RESISTOR T1 T2 PARAMS: RESISTANCE=1k 
R1 T1 T2 {RESISTANCE}
.ends RESISTOR
